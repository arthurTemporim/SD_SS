library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity deslocador_bit is
	port (
	);
end deslocador_bit;

architecture Behavioral of deslocador_bit is

begin


end Behavioral;

