library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity projeto1 is
	port(
		e : in  std_logic_vector (3 downto 0) := "0000"
		s : out std_logic_vector (6 downto 0);
	);
end projeto1;

architecture Behavioral of projeto1 is
begin

s(0) <= e(2) + 

end Behavioral;

