library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity codificador is
end codificador;

architecture Behavioral of codificador is

begin


end Behavioral;

